
// Copyright 2024 Filippo Savi
// Author: Filippo Savi <filssavi@gmail.com>
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
`timescale 10 ns / 1 ns
`include "interfaces.svh"

module fp_add (
    input wire clock,
    axi_stream.slave in_a,
    axi_stream.slave in_b,
    axi_stream.master out
);


    /////////////////////////////////////////
    //         stage 1: scale inputs       //
    /////////////////////////////////////////

    
    /////////////////////////////////////////
    //         stage 2: add mantisse       //
    /////////////////////////////////////////

  
    /////////////////////////////////////////
    //     stage 3: normalize result       //
    /////////////////////////////////////////

  
    /////////////////////////////////////////
    //           stage 4: round            //
    /////////////////////////////////////////

    
  
endmodule
