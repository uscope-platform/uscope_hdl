`timescale 10ns / 1ns

module simple_axi_bram_tb ();


endmodule