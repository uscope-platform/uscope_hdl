`timescale 10ns / 1ns
`include "interfaces.svh"

module simple_axi_bram_tb ();


endmodule