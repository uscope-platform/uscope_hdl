// Copyright 2021 University of Nottingham Ningbo China
// Author: Filippo Savi <filssavi@gmail.com>
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
`timescale 10 ns / 1 ns

module AdcProcessing #(
    parameter DATA_PATH_WIDTH = 16,
    parameter DEST_WIDTH = 8,
    parameter USER_WIDTH = 16,
    DATA_BLOCK_BASE_ADDR = 0,
    FAST_DATA_OFFSET = 0,
    FLTER_TAP_WIDTH = 16,
    DECIMATED = 1,
    DENOISING = 0,
    ENABLE_AVERAGE = 0,
    STICKY_FAULT = 0,
    N_CHANNELS = 4,
    MAX_FILTER_TAPS = 256,
    parameter [N_CHANNELS-1:0] OUTPUT_SIGNED = {N_CHANNELS{1'b1}},
    FILTER_WORKING_WIDTH = DATA_PATH_WIDTH > FLTER_TAP_WIDTH ? DATA_PATH_WIDTH : FLTER_TAP_WIDTH,
    parameter [FLTER_TAP_WIDTH-1:0] FILTER_TAPS [MAX_FILTER_TAPS:0] = '{MAX_FILTER_TAPS+1{0}},
    LINEARIZER_SEGMENTS = 4,
    parameter [DATA_PATH_WIDTH-1:0] LINEARIZER_BOUNDS [N_CHANNELS-1:0][LINEARIZER_SEGMENTS-1:0] = '{default:0},
    parameter [DATA_PATH_WIDTH:0] LINEARIZER_GAINS [N_CHANNELS-1:0][LINEARIZER_SEGMENTS-1:0] = '{default:0},
    PRAGMA_MKFG_MODULE_TOP = "AdcProcessing",
    parameter PRAGMA_MKFG_DATAPOINT_NAMES = "" 
)(
    input  wire       clock,
    input  wire       reset,
    axi_stream.slave  data_in,
    axi_stream.master filtered_data_out,
    axi_stream.master fast_data_out,
    axi_lite.slave    axi_in,
    output reg        fault
);


    initial begin
        $display("--------------------------------------------------------------");
        $display("%s", PRAGMA_MKFG_DATAPOINT_NAMES);
        $display("--------------------------------------------------------------");
    end

    wire shift_enable;
    wire [1:0] latch_mode;
    wire [1:0] clear_latch;
    wire [1:0] trip_high;
    wire [1:0] trip_low;
    wire [7:0] decimation_ratio;

    wire denoise_enable;
    wire signed [DATA_PATH_WIDTH-1:0] denoise_tresh_p [N_CHANNELS-1:0];
    wire signed [DATA_PATH_WIDTH-1:0] denoise_tresh_n [N_CHANNELS-1:0];


    wire signed [DATA_PATH_WIDTH-1:0] comparator_thresholds [0:7];

    wire signed [DATA_PATH_WIDTH-1:0] offset [N_CHANNELS-1:0];
    wire [DATA_PATH_WIDTH-1:0] shift [N_CHANNELS-1:0];

    wire [7:0] n_taps;
    wire [FLTER_TAP_WIDTH-1:0] taps_data;
    wire [7:0] taps_addr;
    wire taps_we, linearizer_enable;

    AdcProcessingControlUnit #(
        .STICKY_FAULT(STICKY_FAULT),
        .DENOISING(DENOISING),
        .FLTER_TAP_WIDTH(FLTER_TAP_WIDTH),
        .DATA_PATH_WIDTH(DATA_PATH_WIDTH),
        .N_CHANNELS(N_CHANNELS)
    ) AdcCU(
        .clock(clock),
        .reset(reset),
        .axi_in(axi_in),
        .data_in_valid(data_in.valid),
        // COMPARATORS
        .comparator_thresholds(comparator_thresholds),
        .latch_mode(latch_mode),
        .clear_latch(clear_latch),
        .trip_high(trip_high),
        .trip_low(trip_low),
        // CALIBRATION
        .shift(shift),
        .offset(offset),
        .shift_enable(shift_enable),
        .fault(fault),
        .linearizer_enable(linearizer_enable),
        // DENOISING
        .denoise_enable(denoise_enable),
        .denoise_tresh_p(denoise_tresh_p),
        .denoise_tresh_n(denoise_tresh_n),
        // FILTERING AND DECIMATION
        .decimation_ratio(decimation_ratio),
        .n_taps(n_taps),
        .taps_data(taps_data),
        .taps_addr(taps_addr),
        .taps_we(taps_we)
    );

    comparator #(
        .DATA_PATH_WIDTH(DATA_PATH_WIDTH)
    )fast_cmp(
        .clock(clock),
        .reset(reset),
        .thresholds(comparator_thresholds[0:3]),
        .data_in(data_in),
        .latching_mode(latch_mode[0]),
        .clear_latch(clear_latch[0]),
        .trip_high(trip_high[0]),
        .trip_low(trip_low[0])
    );

    axi_stream #(
        .DATA_WIDTH(DATA_PATH_WIDTH)
    ) cal_out();

    calibration #(
        .DATA_PATH_WIDTH(DATA_PATH_WIDTH),
        .N_CHANNELS(N_CHANNELS),
        .DATA_BLOCK_BASE_ADDR(DATA_BLOCK_BASE_ADDR),
        .OUTPUT_SIGNED(OUTPUT_SIGNED)
    ) calibrator(
        .clock(clock),
        .reset(reset),
        .data_in(data_in),
        .shift(shift),
        .offset(offset),
        .shift_enable(shift_enable),
        .data_out(cal_out)
    );

    axi_stream #(
        .DATA_WIDTH(DATA_PATH_WIDTH)
    ) denoise_out();

    denoiser #(
        .DATA_PATH_WIDTH(DATA_PATH_WIDTH),
        .DATA_BLOCK_BASE_ADDR(DATA_BLOCK_BASE_ADDR),
        .N_CHANNELS(N_CHANNELS)
    )denoise(
        .clock(clock),
        .reset(reset),
        .thresh_p(denoise_tresh_p),
        .thresh_n(denoise_tresh_n),
        .enable(denoise_enable),
        .data_in(cal_out),
        .data_out(denoise_out)
    );

    axi_stream #(
        .DATA_WIDTH(DATA_PATH_WIDTH)
    ) lin_out();

    linearizer #(
        .DATA_PATH_WIDTH(DATA_PATH_WIDTH),
        .DATA_BLOCK_BASE_ADDR(DATA_BLOCK_BASE_ADDR),
        .N_CHANNELS(N_CHANNELS),
        .DEST_WIDTH(DEST_WIDTH),
        .USER_WIDTH(USER_WIDTH),
        .N_SEGMENTS(LINEARIZER_SEGMENTS),
        .BOUNDS(LINEARIZER_BOUNDS),
        .GAINS(LINEARIZER_GAINS)
    )linearizer(
        .clock(clock),
        .reset(reset),
        .enable(linearizer_enable),
        .data_in(denoise_out),
        .data_out(lin_out)
    );

    assign fast_data_out.data = lin_out.data;
    assign fast_data_out.user = lin_out.user;
    assign fast_data_out.valid = lin_out.valid;
    assign fast_data_out.dest = lin_out.dest + FAST_DATA_OFFSET;
    
    generate
        if(DECIMATED==0)begin
            assign filtered_data_out.data = lin_out.data;
            assign filtered_data_out.valid = lin_out.valid;
            assign filtered_data_out.user = lin_out.user;
            assign filtered_data_out.dest = lin_out.dest;
            assign lin_out.ready = filtered_data_out.ready;

        end else if(DECIMATED==1)begin
            
            standard_decimator #(
                .MAX_DECIMATION_RATIO(16),
                .DATA_WIDTH(DATA_PATH_WIDTH),
                .AVERAGING(ENABLE_AVERAGE),
                .N_CHANNELS(N_CHANNELS)
            ) dec(
                .clock(clock),
                .reset(reset),
                .data_in(lin_out),
                .data_out(filtered_data_out),
                .decimation_ratio(decimation_ratio)
            );

        end else if(DECIMATED == 2)begin


        axi_stream #(
            .DATA_WIDTH(DATA_PATH_WIDTH)
        ) raw_filtered_out();

        fir_filter_serial #(
            .DATA_PATH_WIDTH(DATA_PATH_WIDTH),
            .TAP_WIDTH(FLTER_TAP_WIDTH),
            .MAX_N_TAPS(MAX_FILTER_TAPS),
            .TAPS_IV(FILTER_TAPS)
        )filter(
            .clock(clock),
            .reset(reset),
            .n_taps(n_taps),
            .tap_data(taps_data),
            .tap_addr(taps_addr),
            .tap_write(taps_we),
            .data_in(lin_out),
            .data_out(raw_filtered_out)
        );

        standard_decimator #(
            .MAX_DECIMATION_RATIO(16),
            .DATA_WIDTH(DATA_PATH_WIDTH),
            .AVERAGING(0),
            .N_CHANNELS(N_CHANNELS)
        ) dec(
            .clock(clock),
            .reset(reset),
            .data_in(raw_filtered_out),
            .data_out(filtered_data_out),
            .decimation_ratio(decimation_ratio)
        );
        end
    endgenerate

    axi_stream #(
        .DATA_WIDTH(DATA_PATH_WIDTH)
    ) slow_cmp_in();

    assign slow_cmp_in.data = filtered_data_out.data;
    assign slow_cmp_in.valid = filtered_data_out.valid;
    assign slow_cmp_in.dest = filtered_data_out.dest;

    comparator #(
        .DATA_PATH_WIDTH(DATA_PATH_WIDTH)
    ) slow_cmp(
        .clock(clock),
        .reset(reset),
        .thresholds(comparator_thresholds[4:7]),
        .data_in(slow_cmp_in),
        .latching_mode(latch_mode[1]),
        .clear_latch(clear_latch[1]),
        .trip_high(trip_high[1]),
        .trip_low(trip_low[1])
    );


endmodule
