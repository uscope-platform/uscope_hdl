// Copyright 2024 Filippo Savi
// Author: Filippo Savi <filssavi@gmail.com>
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`timescale 10 ns / 1 ns
`include "interfaces.svh"

module stream_fault_detector #(
    parameter N_CHANNELS = 4,
    parameter STARTING_DEST = 0
)(
    input wire clock,
    input wire reset,
    axi_stream.watcher  data_in,
    axi_lite.slave    axi_in,
    input wire clear_fault,
    output wire        fault
);

    reg [31:0] cu_write_registers [5:0];
    reg [31:0] cu_read_registers  [5:0];


    axil_simple_register_cu #(
        .N_READ_REGISTERS(6),
        .N_WRITE_REGISTERS(6),
        .REGISTERS_WIDTH(32),
        .ADDRESS_MASK('hff)
    ) CU (
        .clock(clock),
        .reset(reset),
        .input_registers(cu_read_registers),
        .output_registers(cu_write_registers),
        .axil(axi_in)
    );


    reg fast_fault = 0;
    reg slow_fault = 0;

    assign fault = fast_fault | slow_fault;

    wire signed [31:0] fast_thresholds [1:0];
    wire signed [31:0] slow_thresholds [1:0];
    wire [7:0] slow_trip_duration;

    assign slow_thresholds[0] = cu_write_registers[0][31:0];
    assign slow_thresholds[1] = cu_write_registers[1][31:0];
    assign slow_trip_duration = cu_write_registers[2][7:0];
    assign fast_thresholds[0] = cu_write_registers[3][31:0];
    assign fast_thresholds[1] = cu_write_registers[4][31:0];

    assign cu_read_registers[4:0] = cu_write_registers[4:0];
    assign cu_read_registers[5] = {fast_fault, slow_fault};


    wire signed[data_in.DATA_WIDTH-1:0] signed_data = $signed(data_in.data);
    wire [7:0] current_address = data_in.dest - STARTING_DEST;

    wire slow_trip = ($signed(signed_data) < $signed(slow_thresholds[0]) || $signed(signed_data) > $signed(slow_thresholds[1])) & ~fast_trip;
    wire fast_trip =  $signed(signed_data) < $signed(fast_thresholds[0]) || $signed(signed_data) > $signed(fast_thresholds[1]);

    reg [7:0] slow_trip_counter [N_CHANNELS-1:0] = '{N_CHANNELS{8'h0}};


    always @(posedge clock) begin
        if(~reset)begin
            fast_fault <= 0;
            slow_fault <= 0;
        end else begin
            if(slow_fault || fast_fault)begin
                if(clear_fault)begin
                    slow_fault <= 0;
                    fast_fault <= 0;
                    slow_trip_counter <= '{N_CHANNELS{8'h0}};
                end
            end else begin
                if(data_in.valid) begin
                    if(fast_trip) begin
                        fast_fault <= 1;
                    end
                    if(slow_trip) begin
                        slow_trip_counter[current_address] <= slow_trip_counter[current_address] + 1;
                    end
                    if(slow_trip_counter[current_address] != 0 & !slow_trip)begin
                        slow_trip_counter[current_address] <= 0;
                    end
                end
                    if(slow_trip_counter[current_address]==slow_trip_duration && slow_trip_duration != 0) begin
                        slow_fault <= 1;
                    end
            end
        end
    end



endmodule


 /**
       {
        "name": "stream_fault_detector",
        "type": "peripheral",
        "registers":[
            {
                "name": "slow_tresh_low",
                "offset": "0x0",
                "description": "Slow fault lower treshold",
                "direction": "RW"
            },
            {
                "name": "slow_tresh_high",
                "offset": "0x4",
                "description": "Slow fault higher treshold",
                "direction": "RW"
            },
            {
                "name": "slow_trip_duration",
                "offset": "0x8",
                "description": "Number of cycles after which a slow fault is triggered",
                "direction": "RW"
            },
            {
                "name": "fast_tresh_low",
                "offset": "0xC",
                "description": "Fast fault lower treshold",
                "direction": "RW"
            },
            {
                "name": "fast_tresh_high",
                "offset": "0x10",
                "description": "Fast fault higher treshold",
                "direction": "RW"
            }
        ]
    }  
    **/
