// Copyright 2021 University of Nottingham Ningbo China
// Author: Filippo Savi <filssavi@gmail.com>
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`timescale 10ns / 1ns
`include "interfaces.svh"
`include "axis_BFM.svh"
							
module register_slice_tb();

    reg  clk, reset;
    axi_stream input_stream();
    axi_stream output_stream();
    //clock generation
    initial clk = 0; 
    always #0.5 clk = ~clk; 
    
    register_slice #(
        .DATA_WIDTH(32),
        .DEST_WIDTH(32),
        .USER_WIDTH(32),
        .N_STAGES(3),
        .READY_REG(0)
    ) UUT(
        .clock(clk),
        .reset(reset),
        .in(input_stream),
        .out(output_stream)
    );


    initial begin
        reset <=1'h1;
        #1 reset <=1'h0;
        output_stream.ready <= 1;
        //TESTS
        #5.5 reset <=1'h1;
        forever begin
            randomize();
            input_stream.user <= $urandom %15;
            input_stream.dest <= $urandom %15;
            input_stream.data <= $urandom;
            input_stream.tlast <= $urandom %2;
            input_stream.valid <= 1;
            #1 input_stream.valid <= 0;
            #10;
        end
    end

endmodule