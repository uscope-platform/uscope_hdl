module fp_fti_tb();


endmodule