// Copyright 2021 University of Nottingham Ningbo China
// Author: Filippo Savi <filssavi@gmail.com>
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`timescale 10 ns / 1 ns

module saturating_adder #(parameter DATA_WIDTH = 32) (
    input wire signed [ DATA_WIDTH-1 :0] a,
    input wire signed [ DATA_WIDTH-1 :0] b,
    input wire signed [ DATA_WIDTH-1 :0] satp,
    input wire signed [ DATA_WIDTH-1 :0] satn,
    output reg signed [ DATA_WIDTH-1 :0] out
);

    reg signed [ DATA_WIDTH :0] int_sum;

    always @(*) begin
        int_sum <= a+b;
        if(int_sum>satp) out <= satp;
        else if(int_sum<satn) out <= satn;
        else out <= int_sum[DATA_WIDTH-1:0];
    end

endmodule