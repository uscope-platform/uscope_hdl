// Copyright 2025 Filippo Savi
// Author: Filippo Savi <filssavi@gmail.com>
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`timescale 10ns / 1ns

module triangle_core #(
    integer N_PARAMETERS = 16,
    integer TIMEBASE_WIDTH = 24
)(
    input wire clock,
    input wire reset,
    input wire trigger,
    input wire [31:0] parameters[N_PARAMETERS-1:0],
    axi_stream.master data_out
);


    wire [31:0] dc_offset;
    assign dc_offset = parameters[0];

    wire [31:0] amplitude;
    assign amplitude = parameters[1];

    wire [31:0] period;
    assign period = parameters[2];

    wire [31:0] phase;
    assign phase = parameters[3];

    wire [31:0] duty;
    assign duty = parameters[4];

    wire [31:0] ramp_increment;
    assign ramp_increment = parameters[5];

    wire [31:0] dest_out;
    assign dest_out = parameters[6];

    wire [31:0] user_out;
    assign user_out = parameters[7];


    reg[TIMEBASE_WIDTH-1:0] generator_counter = 0;
    reg running = 0;

    initial begin
        data_out.data = 0;
        data_out.dest = 0;
        data_out.tlast = 0;
        data_out.valid = 0;
        data_out.user = 0;
    end


    wire down_ramp;
    assign down_ramp = generator_counter > duty-1;

    always_ff@(posedge clock)begin
        data_out.tlast <= 0;
        data_out.valid <= 0;
        if(!running)begin
            if(trigger)begin
                running <= 1;
            end
            generator_counter <= phase;
        end else begin
            if(trigger)begin
                if(generator_counter==period-1)begin
                    generator_counter <= 0;
                end else begin
                    if(down_ramp) begin
                        generator_counter <= generator_counter-ramp_increment;
                    end else begin
                        generator_counter <= generator_counter+ramp_increment;
                    end
                end
                data_out.data <= generator_counter;
                data_out.dest <= dest_out;
                data_out.user <= user_out;
                data_out.valid <= 1;
                data_out.tlast <= 1;

            end
        end
    end


    always_comb begin

    end

endmodule
